module SUB44(
	input logic signed [3:0] A, B, 
	output logic signed [4:0] D); 

	  assign D = A-B ;
endmodule

