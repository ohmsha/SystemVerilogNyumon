module parameter_update(input logic [31:0] IN, output logic [31:0] OUT);
   defparam I0.PARAM=10'd256;
   parameter_example  I0  (.*);
endmodule // parameter_update
