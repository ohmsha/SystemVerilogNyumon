module SUB4(
	input logic [3:0] A, B, 
	output logic [3:0] D); 

	  assign D = A-B ;
endmodule

