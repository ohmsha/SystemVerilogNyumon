module parameter_update(input logic [31:0] IN, output logic [31:0] OUT);
   parameter_example  #(.PARAM(10'd256)) I0  (.*);
endmodule // parameter_update

